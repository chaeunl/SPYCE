.param w_0_0_0=1.2257267517233448 w_0_0_1=0.4986420275972627 w_0_0_2=1.77809112619885 w_0_0_3=1.536309053688945 w_0_1_0=1.4844877122006945 w_0_1_1=0.9279773441646544 w_0_1_2=-0.9519885422026324 w_0_1_3=0.5047848031780162 w_0_2_0=0.23809536877768012 w_0_2_1=1.6258771187692593 w_0_2_2=-0.8232887181810853 w_0_2_3=2.1825927902884823 w_1_0_0=0.8759648247704082 w_1_0_1=-0.532554904948053 w_1_0_2=2.1612867771304614 w_1_0_3=1.4346993699716757 w_1_1_0=1.450491332504237 w_1_1_1=1.7349468046489727 w_1_1_2=0.38089822075805935 w_1_1_3=0.14117991030025712 w_1_2_0=0.45933913372199386 w_1_2_1=0.022378765256725552 w_1_2_2=1.022235370297886 w_1_2_3=-0.18468851747648873 
.param a_0_0_0=1.1053176424612605 a_0_0_1=0.5707876204821543 a_0_0_2=1.8606583931178133 a_0_0_3=1.4846270963462818 a_0_1_0=-0.5054963630374931 a_0_1_1=1.2574519309663121 a_0_1_2=0.547825027306895 a_0_1_3=-0.11890338356953922 a_0_2_0=-0.4798406358519117 a_0_2_1=-0.5454931594832195 a_0_2_2=1.3379475198595174 a_0_2_3=0.005937917602876652 a_1_0_0=-0.8026606115286551 a_1_0_1=1.2037933590150134 a_1_0_2=-0.40003885907593606 a_1_0_3=1.3584496589718436 a_1_1_0=1.620875159013401 a_1_1_1=1.1978907551923323 a_1_1_2=0.9379324281508752 a_1_1_3=1.1882424712948518 a_1_2_0=1.3125428606476404 a_1_2_1=0.804157891312165 a_1_2_2=0.9398795495705174 a_1_2_3=1.4644389807004243 
.param vt_0_0_0=0.3832479167757694 vt_0_0_1=1.0181219284303653 vt_0_0_2=1.4342456018596295 vt_0_0_3=1.1966667793893717 vt_0_1_0=1.056378770001463 vt_0_1_1=1.4525463606007811 vt_0_1_2=2.1500313236358974 vt_0_1_3=1.7049333577948378 vt_0_2_0=0.43225609558752276 vt_0_2_1=0.42728926935327305 vt_0_2_2=1.4695535494690977 vt_0_2_3=0.11503096456236683 vt_1_0_0=1.1955018379931541 vt_1_0_1=1.6404962459905894 vt_1_0_2=-0.05045473349032892 vt_1_0_3=0.04818882945205205 vt_1_1_0=0.18705942711884394 vt_1_1_1=2.1011753648091602 vt_1_1_2=-0.15466181714360827 vt_1_1_3=-0.3308210964579007 vt_1_2_0=2.2202164590276716 vt_1_2_1=0.015803976783475004 vt_1_2_2=-0.7536113706161204 vt_1_2_3=1.4312221945842754 
* open file
